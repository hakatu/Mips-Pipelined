library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity instruction_memory is
    Port ( address : in  STD_LOGIC_VECTOR (31 downto 0);
           clk: in STD_logic;
           Instr : out  STD_LOGIC_VECTOR (31 downto 0));
end entity;


architecture behavioral of instruction_memory is

type ARRAY_256 is ARRAY (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
--hexcode trong
--signal MemContent: ARRAY_256 := (   X"0c000004",
--X"20090001",
--X"ac090000",
--X"15200002",
--X"200a0002",
--X"03e00008",
--X"08000008",
--X"200b0003",
--X"a00a0001",
--X"8c0c0000",
--X"800d0001",
--X"20090005",
--X"21280000",
--X"200a0000",
--X"200b0000",
--X"200cffff",
--X"200d0000",
--X"200e0000",
--X"200f0000",
--X"012c4820",
--X"012c5020",
--X"01005820",
--X"11200004",
--X"1140fffb",
--X"010b4020",
--X"014c5020",
--X"08000017",
--X"ac080004",
--X"20090000",
--X"20080000",
--X"200a0000",
--X"200b0000",
--X"200c0000",
--X"200d0000",
--X"200e0000",
--X"200f0000",
--X"20100002",
--X"02108820",
--X"02319020",
--X"02529820",
--X"0273a020",
--X"0294a820",
--X"02b5b020",
--X"02d6b820",
--X"02f74020",
--X"01084820",
--X"01295020",
--X"014a5820",
--X"016b6020",
--X"018c6820",
--X"01ad7020",
--X"01ce7820",
--X"01efc020",
--X"0318c820",
--X"03392020",
--X"00842820",
--X"00a53020",
--X"00c63820",
--X"00e71020",
--X"00421820",
--X"ac030014",
--X"20090000",
--X"20080000",
--X"200a0000",
--X"200b0000",
--X"200c0000",
--X"200d0000",
--X"200e0000",
--X"200f0000",
--X"20080002",
--X"1208001b",
--X"02108820",
--X"02319020",
--X"02529820",
--X"0273a020",
--X"0294a820",
--X"02b5b020",
--X"02d6b820",
--X"0800005f",
--X"02f74020",
--X"01084820",
--X"01295020",
--X"014a5820",
--X"016b6020",
--X"018c6820",
--X"01ad7020",
--X"01ce7820",
--X"01efc020",
--X"0318c820",
--X"08000045",
--X"03392020",
--X"00842820",
--X"00a53020",
--X"00c63820",
--X"08000045",
--X"00e71020",
--X"00421820",
--X"0800005a",
--X"ac170024",
--X"00000000",--0 toi 144
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--154 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--164 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--184 20 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--204 20 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--224 20 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--244 20 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--254 10 dong
--X"00000000", --211
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--221 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--231 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--241 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",--251 10 dong
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000",
--X"00000000"
--);

signal MemContent: ARRAY_256 := (   X"20090005",X"21280000",X"200a0000",X"200b0000",X"200cffff",X"200d0000",X"200e0000",X"200f0000",X"012c4820",X"012c5020",X"01005820",X"11200004",X"1140fffb",X"010b4020",X"014c5020",X"0800000c",X"ac080004",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000" );
--hex code test jump 
--signal MemContent: ARRAY_256 := (   X"200b0003",X"ac0b0000",X"8c0a0000",X"116a0001",X"014b4820",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000" );
----hex code checkloi
--signal MemContent: ARRAY_256 :=	(	X"20090001",X"200a0001",X"200b0000",X"ad690000",X"216b0004",X"ad6a0000",X"216b0004",X"20080000",X"012a6020",X"000a4820",X"000c5020",X"ad6c0000",X"216b0004",X"21080001",X"2001000f",X"1428fff8",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--											X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"	);
----hex code fibonacci(thieu sub)
--signal MemContent: ARRAY_256 := (   X"0c000002",X"01e00008",X"20090001",X"31290003",X"35290003",X"200a0001",X"012a5824",X"012a6025",X"012a6827",X"00094842",X"000a5040",X"112a0003",X"200f0005",X"152a0002",X"200f0004",X"012a702a",X"292e000a",
--                                            X"ac090000",X"8c0a0000",X"a009000a",X"800a000a",X"200f0064",X"08000001",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000" );
--testcodefinal
--signal MemContent: ARRAY_256 := (   X"0c000002",X"ac1f0000",X"21290001",X"21ef0001",X"01bf6820",X"03e00008",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000" );
-----testcode jr va jal
--signal MemContent: ARRAY_256 := (   X"200d4e20",X"ac0d0008",X"8c0d0008",X"a00d0013",X"800f0013",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000" );
-----test sb lb lw sw
--signal MemContent: ARRAY_256 := ( "10010000000111100000000000110010",
--"00100011110111100000000000000001",
--"00100000000000010000000000000001",
--"00100000000001010000000000000000",
--"00010000001111100000000000000011",
--"00000000101000010010100000100000",
--"00100000001000010000000000000001",
--"00001000000000000000000000000100",
--"00100000000000010000000000000001",
--"00100000000001100000000000000000",
--"00010000001111100000000000000101",
--"00000000001000000001000000100000",
--"00000000001000000001100000100000",
--"00001100000000000000000001101111",
--"00000000110001000011000000100000",
--"00001000000000000000000000001010",
--"00100000000000010000000000000011",
--"00100000000000100000000000000001",
--"00100000000000110000000000000001",
--"00010000001111100000000000000101",
--"00000000010000110010000000100000",
--"00100000011000100000000000000000",
--"00100000100000110000000000000000",
--"00100000001000010000000000000001",
--"00001000000000000000000000010011",
--"00100000011001110000000000000000",
--"00100000000000010000000000000000",
--"00100000000000110000000000000001",
--"00010000001111100000000000000101",
--"00100000001000100000000000000001",
--"00001100000000000000000001101111",
--"00100000100000110000000000000000",
--"00100000001000010000000000000000",
--"00001000000000000000000000011100",
--"00100000011010000000000000000000",
--"00100000000000010000000000000001",
--"10001100000111100000000000110010",
--"00100000000000100000000000100001",
--"00010000001000100000000000001000",
--"00110011110001000000000000000001",
--"00010100100000000000000000000010",
--"00100001010010100000000000000001",
--"00001000000000000000000000101100",
--"00100001001010010000000000000001",
--"00100000001000010000000000000001",
--"00000000000111101111000001000010",
--"00001000000000000000000000100110",
--"10010000000010110000000000000001",
--"10010000000011000000000000000010",
--"10010000000011010000000000000011",
--"10010000000011100000000000000100",
--"10010000000011110000000000000101",
--"10010000000100000000000000000110",
--"10010000000100010000000000000111",
--"10010000000100100000000000001000",
--"10010000000100110000000000001001",
--"00100000000000010000000000000001",
--"00100000000001000000000000001010",
--"00010000001001000000000000101010",
--"00100001011000100000000000000000",
--"00100001100000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010010110000000000000000",
--"00100000011011000000000000000000",
--"00100001100000100000000000000000",
--"00100001101000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010011000000000000000000",
--"00100000011011010000000000000000",
--"00100001101000100000000000000000",
--"00100001110000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010011010000000000000000",
--"00100000011011100000000000000000",
--"00100001110000100000000000000000",
--"00100001111000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010011100000000000000000",
--"00100000011011110000000000000000",
--"00100001111000100000000000000000",
--"00100010000000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010011110000000000000000",
--"00100000011100000000000000000000",
--"00100010000000100000000000000000",
--"00100010001000110000000000000000",
--"00001100000000000000000001110111",
--"00100000010100000000000000000000",
--"10101100000111010000000000101100"
--);
--signal MemContent: ARRAY_256 := (   X"200f000d",X"ac0f0014",X"8c080014",X"20090001",X"00005020",X"200d0001",X"01205820",X"012a4820",X"01605020",X"0128602a",X"118dfffb",X"11280002",X"200d0037",X"0800000f",X"200d0064",X"ac0d0018",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
--                            X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000");
begin
Instr <= MemContent(to_integer(unsigned(address(31 downto 2))));
end behavioral;